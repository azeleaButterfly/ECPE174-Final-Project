module rng_testbench ();
    


    initial begin
        
    end
endmodule