module simon_says(
    
);


endmodule